module pattern2(row_bin, col);
	input [3:0]	row_bin;
	output	reg [15:0]	col;
	
	// 小綠人行走圖形編碼2
	// 紅色為1 黃色為0
	always@ (*) begin
		case (row_bin)
			4'd0:	col=16'b0000000000000000;
			4'd1:	col=16'b0000110000000000;
			4'd2:	col=16'b0001111000000000;
			4'd3:	col=16'b0000110000000000;
			4'd4:	col=16'b0000011000000000;
			4'd5:	col=16'b0000011100000000;
			4'd6:	col=16'b0000011010000000;
			4'd7:	col=16'b0000011110000000;
			4'd8:	col=16'b0000001110000000;
			4'd9:	col=16'b0000001100000000;
			4'd10:	col=16'b0000001100000000;
			4'd11:	col=16'b0000011100000000;
			4'd12:	col=16'b0000010010000000;
			4'd13:	col=16'b0000001001000000;
			4'd14:	col=16'b0000111000100000;
			4'd15:	col=16'b0000000000000000;
			default:col=16'b0000000000000000;
		endcase
	end
endmodule